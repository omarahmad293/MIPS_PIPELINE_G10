module Shiftleft2_32(IN,Out);
input[31:0] IN;
output[31:0] Out;

assign Out = IN<<2;


endmodule
